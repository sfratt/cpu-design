library ieee;
use ieee.std_logic_1164.all;

entity d_cache is
    port(

    );
end d_cache;

architecture d_cache_arch of d_cache is

    signal 

begin

end architecture d_cache_arch;