library ieee;
use ieee.std_logic_1164.all;

entity data_cache is
    port(

    );
end data_cache;

architecture d_cache_arch of data_cache is

    signal 

begin

end architecture d_cache_arch;